* MAX4224 CLOSED LOOP GAIN RESPONSE GAIN = +2
* 4224AVCL.CIR
*NOTE OFFSET OF AMPLIFIER MUST BE ZERO !
*
*  
XAR1 3 2 7 4 6 MAX4224
*   +IN -IN VCC VEE OUT             
VP 7 0  5V
VN 4 0  -5V
VIN 3 0 AC 1
RF 6 2 470
RG 2 0 470
RL 6 0 100
.OPTIONS RELTOL=.01
.AC DEC 10 1 10000meg               
.PROBE                             
.LIB MAX4223.FAM
.END


