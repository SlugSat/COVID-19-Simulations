* OPA855 - Rev. A
* Created by Sean Cashin; December 16, 2019
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2019 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT OFFSET VOLTAGE VS. TEMPERATURE (Vos Drift)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt OPA855 IN+ IN- VCC VEE OUT
******************************************************
.MODEL              R_NOISELESS RES (T_ABS=-273.15)
***                 
C_C1                MID CLAMP 20p
C_C1a               N1492098 N1492108 19.9p
C_C1a1              MID N1492376 4f
C_C1a15             N1483677 N1483687 29.36p
C_C1a16             PSRRP N1481259 50p
C_C1a17             N1483713 PSRRN 34.6f
C_C1a35             N1461236 N1461246 18.72p
C_C1a36             N1461252 CMRR 53f
C_C1a39             N1481243 N1481253 22.74p
C_C1a40             N1483693 N1483703 34.6f
C_C33               N406634 0 1e-15
C_C34               N317950 0 1
C_C35               N406794 0 1e-15
C_C44               N1446217 MID 3p
C_C46               N1507810 N1508339 5.3f
C_C7                N31014 MID 1p
C_C8                MID N35813 1e-15
C_C9                MID N38096 1e-15
C_C_CMn             MID ESDN 0.6p
C_C_CMn1            ESDN ESDP 0.2p
C_C_CMp             ESDP MID 0.6p
C_C_VIMON           MID VIMON 1e-12
C_C_VOUT_S          MID VOUT_S 1e-12
E_E3                N112292 MID OUT MID 1
E_E6                MID 0 N317950 0 1
G_G1                N1492098 MID N1446217 ZO -1.75
G_G111              N1461252 MID N1461246 MID 333
G_G114              N1481243 MID VCC_B MID 0.716
G_G115              N1481259 MID N1481253 MID 4
G_G116              N1483677 MID VEE_B MID 1.578
G_G12               N1446199 MID N1507810 MID -1
G_G2                N10570 N10561 CMRR MID -1e-3
G_G36               VCC_B 0 VCC 0 -1
G_G37               VEE_B 0 VEE 0 -1
G_G4                N1254860 MID N1492126 MID -130
G_G5                N1492118 MID N1492108 MID -1
G_G6                N25816 N11984 PSRRP PSRRN -1e-3
G_G76               N1461236 MID ESDP MID 117m
G_G77               N1483693 MID N1483687 MID 21.74
G_G78               N1483713 MID N1483703 MID 21.74
G_G8                VCC_CLP MID N35813 MID -1E-3
G_G9                VEE_CLP MID N38096 MID -1E-3
G_G95               N1508339 MID CLAMP MID -3.5
I_I_B               N06456 MID DC 12u
I_I_OS              ESDN MID DC 12.1u
I_I_Q               VCC VEE DC 16.4m
L_L1                N1446199 N1446217 200p
L_L2                PSRRP N1490067 4n
R_R1                ESDP IN+ R_NOISELESS 10e-3
R_R10               ESDN N11991 R_NOISELESS 1e-3
R_R107              VCC_B 0 R_NOISELESS 1
R_R108              N317950 0 R_NOISELESS 1e12
R_R109              VEE_B 0 R_NOISELESS 1
R_R110              VCC_B N406634 R_NOISELESS 1e-3
R_R111              N406634 N317950 R_NOISELESS 1e6
R_R112              N317950 N406794 R_NOISELESS 1e6
R_R113              N406794 VEE_B R_NOISELESS 1e-3
R_R146              N1461236 MID R_NOISELESS 1
R_R147              N1461252 MID R_NOISELESS 1
R_R148              N1483713 MID R_NOISELESS 1
R_R162              ESDN ESDP R_NOISELESS 5k
R_R1a               N1492108 N1492098 R_NOISELESS 10e3
R_R1a1              N1492126 N1492118 R_NOISELESS 14k
R_R1a14             N1461236 N1461246 R_NOISELESS 10e3
R_R1a15             N1461252 CMRR R_NOISELESS 10e3
R_R1a16             PSRRP MID R_NOISELESS 2.8
R_R1a17             N1483693 N1483703 R_NOISELESS 10e3
R_R1a18             N1483713 PSRRN R_NOISELESS 10e3
R_R1a40             N1481243 N1481253 R_NOISELESS 10e3
R_R1a41             N1490067 N1481259 R_NOISELESS 7
R_R1a42             N1483677 N1483687 R_NOISELESS 10e3
R_R2                ESDN IN- R_NOISELESS 10e-3
R_R21               N11984 N25816 R_NOISELESS 1e3
R_R211              MID N1254860 R_NOISELESS 1
R_R225              MID N1446199 R_NOISELESS 1
R_R226              MID N1446217 R_NOISELESS 35
R_R227              N1508339 MID R_NOISELESS 1
R_R228              N1507810 MID R_NOISELESS 4.28k
R_R229              N1508339 N1507810 R_NOISELESS 10k
R_R241              MID CLAMP R_NOISELESS 6.4k
R_R245              VCC VEE R_NOISELESS 4.5k
R_R246              N1481243 MID R_NOISELESS 1
R_R247              N1481259 MID R_NOISELESS 1
R_R248              N1483677 MID R_NOISELESS 1
R_R249              N1483693 MID R_NOISELESS 1
R_R25               MID N28602 R_NOISELESS 1e9
R_R250              MID N1492098 R_NOISELESS 1
R_R26               N30136 MID R_NOISELESS 1e9
R_R27               MID N30913 R_NOISELESS 1
R_R28               N31014 N30913 R_NOISELESS 1e-3
R_R29               N35675 VCC_B R_NOISELESS 1e3
R_R2a               MID N1492108 R_NOISELESS 13.33k
R_R2a1              N1492376 N1492126 R_NOISELESS 10k
R_R2a16             N1483687 MID R_NOISELESS 0.542
R_R2a17             N1483703 MID R_NOISELESS 482.2
R_R2a18             PSRRN MID R_NOISELESS 482.2
R_R2a36             N1461246 MID R_NOISELESS 0.85
R_R2a37             CMRR MID R_NOISELESS 30.1
R_R2a40             N1481253 MID R_NOISELESS 0.7
R_R3                MID ESDP R_NOISELESS 2.3MEG
R_R30               N35813 N35675 R_NOISELESS 1e-3
R_R31               VCC_CLP MID R_NOISELESS 1e3
R_R32               N38050 VEE_B R_NOISELESS 1e3
R_R33               N38096 N38050 R_NOISELESS 1e-3
R_R34               VEE_CLP MID R_NOISELESS 1e3
R_R4                ESDN MID R_NOISELESS 2.3MEG
R_R6                MID N1492118 R_NOISELESS 1
R_R60               MID AOL_1 R_NOISELESS 1
R_R8                N10561 N10570 R_NOISELESS 1e3
R_R81               MID N110431 R_NOISELESS 1e9
R_R83               MID N112292 R_NOISELESS 1e9
R_R9                N10570 N11984 R_NOISELESS 1e-3
R_R_VIMON           VIMON N110431 R_NOISELESS 100
R_R_VOUT_S          VOUT_S N112292 R_NOISELESS 100
R_Rdummy            MID ZO R_NOISELESS 200
R_Rx                ZO N1254860 R_NOISELESS 2k
V_VCM_MAX           N30136 VCC_B -0.4
V_VCM_MIN           N28602 VEE_B 1.1
X_e_n               ESDP N06456 VNSE
X_ESD_OUT           OUT VCC VEE ESD_OUT
X_H3                OUT ZO N110431 MID 08_Op_Amp_Complete_H3
X_i_np1             ESDN MID FEMT
X_IQ_N              MID VIMON MID VEE IQ_SRC
X_IQ_P              VIMON MID VCC MID IQ_SRC
X_U1                MID N06456 FEMT
X_U2                N31014 N11991 AOL_1 MID AOL_1
X_U3                AOL_1 MID CLAMP MID AOL_2
X_U5                VIMON MID N35675 VCC_B CLAWP
X_U6                VIMON MID VEE_B N38050 CLAWN
X_VCM_CLAMP         N25816 MID N30913 MID N30136 N28602 VCM_CLAMP
X_VOS_DRIFT         N749288 N06456 VOS_DRIFT
X_VOS_VS_VCM        N10561 N749288 VCC VEE VOS_VS_VCM
.ENDS OPA855

.subckt 08_Op_Amp_Complete_H3 1 2 3 4  
H_H3         3 4 VH_H3 -1e3
VH_H3         1 2 0V
.ends 08_Op_Amp_Complete_H3

*
.subckt AOL_1 VC+ VC- IOUT+ IOUT-
.param Gain = 1
.param Ipos = .5
.param Ineg = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(Gain*V(VC+,VC-),Ineg,Ipos)}
.ends
*$
*
.subckt AOL_2 VC+ VC- IOUT+ IOUT-
.param Gain = 1
.param Ipos = 0.055
.param Ineg = -0.055
G1 IOUT+ IOUT- VALUE={LIMIT(Gain*V(VC+,VC-),Ineg,Ipos)}
.ends
*$
*
.subckt CLAWn VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {abs(V(VC+,VC-))} =
+(0, 1.02e-3)
+(20.5, 1.19e-3)
+(46.37, 1.37e-3)
+(55.32, 1.43e-3)
+(61.86, 1.47e-3)
+(67.19, 1.51e-3)
+(72.22, 1.55e-3)
+(78.37, 1.60e-3)
+(85.63, 1.63e-3)
+(90.22, 1.67e-3)
+(93.85, 1.70e-3)
+(97.87, 1.74e-3)
+(101.1, 1.76e-3)
+(104.5, 1.80e-3)
+(106.9, 1.83e-3)
+(109.9, 1.91e-3)
+(111.9, 2.026e-3)

.ends
*$
*
.subckt CLAWp VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {abs(V(VC+,VC-))} =
+(0, 7.88e-4)
+(6.1, 8.68e-4)
+(15.2, 9.53e-4)
+(27.1, 1.04e-3)
+(42.8, 1.16e-3)
+(60.7, 1.29e-3)
+(97.11, 1.66e-3)
+(106.7, 1.81e-3)
+(112.2, 1.99e-3)
+(120.1, 2.40e-3)

.ends
*$
*
.subckt ESD_OUT OUT VCC VEE
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=500e-3 Voff=450e-3)
S1 VCC OUT OUT VCC ESD_SW
S2 OUT VEE VEE OUT ESD_SW
.ends
*$
*
.subckt FEMT 1 2
.param FLWF=1000
.param NLFF=33
.param NVRF=2.5
.param GLFF={PWR(FLWF,0.25)*NLFF/1164}
.param RNVF={1.184*PWR(NVRF,2)}
.model DNVF D KF={PWR(FLWF,0.5)/1e11} IS=1.0e-16
I1 0 7 10e-3
I2 0 8 10e-3
D1 7 0 DNVF
D2 8 0 DNVF
E1 3 6 7 8 {GLFF}
R1 3 0 1e9
R2 3 0 1e9
R3 3 6 1e9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1e9
R7 4 0 1e9
G1 1 2 3 4 1e-6
.ends
*$
*
.subckt IQ_SRC VC+ VC- IOUT+ IOUT-
.param Gain = 1e-3
G1 IOUT+ IOUT- VALUE={IF( (V(VC+,VC-)<=0),0,Gain*V(VC+,VC-) )}
.ends
*$
*
.subckt VCM_CLAMP VIN+ VIN- IOUT- IOUT+ VP+ VP-
.param Gain = 1
G1 IOUT+ IOUT- VALUE={LIMIT(Gain*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ends
*$
*
.subckt VNSE 1 2
.param FLW=1000
.param NLF=3
.param NVR=0.98
.param GLF={PWR(FLW,0.25)*NLF/1164}
.param RNV={1.184*PWR(NVR,2)}
.model DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
* Circuit connections
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ends
*$
*
.subckt VOS_DRIFT VOS+ VOS-
.param DC = -4e-4
.param POL = 1
.param DRIFT = 20e-6
E1 VOS+ VOS- VALUE={DC+POL*DRIFT*(TEMP-27)}
.ends
*$
*
.subckt VOS_VS_VCM V+ V- REF+ REF-
* Positive rail Vos
E1 V+ 1 TABLE {(V(REF+, V-))} =
+(0.35, 450e-6)
+(0.4, 435e-6)
+(0.55, 275e-6)
+(0.65, 150e-6)
+(0.75, 75e-6)
+(0.85, 25e-6)
+(1, 0)
* Negative rail Vos
V1 1 V- 0
.ends
*$
*
*$
